// ----------------------------------------
// ----------------------------------------
// Top module for StarSoC game design
// top.sv
// Justin Coppola
// 04/22/2025
// ----------------------------------------
// ----------------------------------------

module top (
    input clk,
    input left_button,
    input right_button,
    input shoot_button,
    output x,
    output y
);

endmodule